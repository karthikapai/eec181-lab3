`timecale 1us / 1us
module lab2(
//FPGA Pins
//Clock Pins
CLOCK_50,
DRAM_CLK,

//SEVEN Segment Display
HEX0,
HEX1,
HEX2,
HEX3,
HEX4,
HEX5,

//Pushbuttons
KEY,

//LEDs
LEDR,

//Slider Switches
//SW,

//HPS Pins
//DDR3 SDRAM
HPS_DDR3_ADDR,
HPS_DDR3_BA,
HPS_DDR3_CAS_N,
HPS_DDR3_CKE,
HPS_DDR3_CK_N,
HPS_DDR3_CK,
HPS_DDR3_CS_N,
HPS_DDR3_DM,
HPS_DDR3_DQ,
HPS_DDR3_DQS_N,
HPS_DDR3_DQS,
HPS_DDR3_ODT,
HPS_DDR3_RAS_N,
HPS_DDR3_RESET_N,
HPS_DDR3_RZQ,
HPS_DDR3_WE_N,
DRAM_ADDR,      // add sdram ports here      
DRAM_BA,        
DRAM_CAS_N,   
DRAM_CKE,       
DRAM_CS_N,    
DRAM_DQ,        
DRAM_UDQM, DRAM_LDQM,       
DRAM_RAS_N,    
DRAM_WE_N
);

//Port Declaration
//FPGA Pins
input CLOCK_50;
output DRAM_CLK;
output [0:6] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
input [3:0] KEY;
output [9:0] LEDR;
//input [9:0] SW;

//HPS Pins
//DDR3 SDRAM
output[14:0] HPS_DDR3_ADDR;  //FIXME: should me 13 bits
output [2:0] HPS_DDR3_BA;
output HPS_DDR3_CAS_N;
output HPS_DDR3_CKE;
output HPS_DDR3_CK_N;
output HPS_DDR3_CK;
output HPS_DDR3_CS_N;
output [3:0] HPS_DDR3_DM;
inout [31:0] HPS_DDR3_DQ;
inout [3:0] HPS_DDR3_DQS_N;
inout [3:0] HPS_DDR3_DQS;
output HPS_DDR3_ODT;
output HPS_DDR3_RAS_N;
output HPS_DDR3_RESET_N;
input HPS_DDR3_RZQ;
output HPS_DDR3_WE_N;

//SDRAM pins
output [12:0] DRAM_ADDR;       
output [1:0]  DRAM_BA;         
output        DRAM_CAS_N;      
output        DRAM_CKE;         
output        DRAM_CS_N;      
inout  [15:0] DRAM_DQ;         
output        DRAM_UDQM, DRAM_LDQM;        
output        DRAM_RAS_N;     
output        DRAM_WE_N;   

//REG/WIRE declarations
wire [31:0] hex5_0bus;
wire [31:0] thirty2bit_in;
wire [31:0] Hex0_Hex5; 

parameter H = 7'b1001000;
parameter E = 7'b0110000;
parameter L = 7'b1110001;
parameter O = 7'b0000001;
parameter U = 7'b1000001;
parameter R = 7'b1111010;
parameter D = 7'b1000010;
parameter space = 7'b1111111;
wire reg [0:11] Helloworld = {H,E,L,L,O,space,U,U,O,R,L,D};
unsigned int i = 0;

int speed = 1000;
wire reg [0:6] hex5, hex4, hex3, hex2, hex1 ,hex0;
assign HEX5 = hex5;
assign HEX4 = hex4;
assign HEX3 = hex3;
assign HEX2 = hex2;
assign HEX1 = hex1;
assign HEX0 = hex0;

always @ (KEY[0] ==1)
begin
# speed;
hex5 = helloworld[(i)%12];
hex4 = helloworld[(i+1)%12];
hex3 = helloworld[(i+2)%12];
hex2 = helloworld[(i+3)%12];
hex1 = helloworld[(i+4)%12];
hex0 = helloworld[(i+5)%12];
i = (i+1) % 12;
if(KEY[1] = 1) begin
speed = speed - 10;
end 
else if begin









//EVERYTHING BELOW HERE WAS (mostly) GENERATED BY QSYS
//Structural Coding


    mysystem u0 (
        .system_ref_clk_clk     (CLOCK_50),                                           //   system_ref_clk.clk
        .system_ref_reset_reset (~KEY[0]),                                               // system_ref_reset.reset
        .to_hex_to_led_export   (thirty2bit_in),    //    to_hex_to_led.export
        .sdram_clk_clk          (DRAM_CLK),                                           //        sdram_clk.clk
        .pushbutton_export      (~KEY[3:1]),                                          //       pushbutton.export
        .hex5_0bus_export       (hex5_0bus),                                          //        hex5_0bus.export
		  //.rled_export            (led),                         //             rled.export
        .memory_mem_a           (HPS_DDR3_ADDR),                                      //           memory.mem_a
        .memory_mem_ba          (HPS_DDR3_BA),          //                 .mem_ba
        .memory_mem_ck          (HPS_DDR3_CK),          //                 .mem_ck
        .memory_mem_ck_n        (HPS_DDR3_CK_N),        //                 .mem_ck_n
        .memory_mem_cke         (HPS_DDR3_CKE),         //                 .mem_cke
        .memory_mem_cs_n        (HPS_DDR3_CS_N),        //                 .mem_cs_n
        .memory_mem_ras_n       (HPS_DDR3_RAS_N),       //                 .mem_ras_n
        .memory_mem_cas_n       (HPS_DDR3_CAS_N),       //                 .mem_cas_n
        .memory_mem_we_n        (HPS_DDR3_WE_N),        //                 .mem_we_n
        .memory_mem_reset_n     (HPS_DDR3_RESET_N),     //                 .mem_reset_n
        .memory_mem_dq          (HPS_DDR3_DQ),          //                 .mem_dq
        .memory_mem_dqs         (HPS_DDR3_DQS),         //                 .mem_dqs
        .memory_mem_dqs_n       (HPS_DDR3_DQS_N),       //                 .mem_dqs_n
        .memory_mem_odt         (HPS_DDR3_ODT),         //                 .mem_odt
        .memory_mem_dm          (HPS_DDR3_DM),          //                 .mem_dm
        .memory_oct_rzqin       (HPS_DDR3_RZQ),         //                 .oct_rzqin
		.sdram_wire_addr        (DRAM_ADDR),        //       sdram_wire.addr
        .sdram_wire_ba          (DRAM_BA),          //                 .ba
        .sdram_wire_cas_n       (DRAM_CAS_N),       //                 .cas_n
        .sdram_wire_cke         (DRAM_CKE),         //                 .cke
        .sdram_wire_cs_n        (DRAM_CS_N),        //                 .cs_n
        .sdram_wire_dq          (DRAM_DQ),          //                 .dq
        .sdram_wire_dqm         ({DRAM_UDQM, DRAM_LDQM}),         //                 .dqm
        .sdram_wire_ras_n       (DRAM_RAS_N),       //                 .ras_n
        .sdram_wire_we_n        (DRAM_WE_N)         //                 .we_n
		  
    );

	        
	 
endmodule


