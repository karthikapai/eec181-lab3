module to_led (
input input_bit,
output led
);

assign led = input_bit;

endmodule
